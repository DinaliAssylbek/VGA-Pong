module glyph_rom(

	// Input signals
	input [5:0] char_index,   // 6-bit character index to select the glyph
	input [2:0] glyph_column, // 3-bit column index within the 8x8 glyph grid
	input [2:0] glyph_row,    // 3-bit row index within the 8x8 glyph grid
	
	// Output signal
	output wire pixel         // Pixel value at the specified row and column for the glyph
	
);
	reg [63:0] glyph; // Register to store the 8x8 glyph as a 64-bit binary value
	
	// Always block to assign the glyph value based on the character index
	always @(*)
		case(char_index)
			// Character Glyphs
			0: glyph = 64'b00000010_00000010_00000010_00011110_00100010_00100010_00011110_00000000;  // P
			1: glyph = 64'b00100010_00010010_00001010_00011110_00100010_00100010_00011110_00000000;  // R
			2: glyph = 64'b00111110_00000010_00000010_00111110_00000010_00000010_00111110_00000000;  // E
			3: glyph = 64'b00011100_00100010_00100000_00011100_00000010_00100010_00011100_00000000;  // S
			4: glyph = 64'b00100010_00100010_00100010_00111110_00100010_00100010_00011100_00000000;  // A
			5: glyph = 64'b00001000_00001000_00001000_00001000_00001000_00001000_00111110_00000000;  // T
			6: glyph = 64'b00011100_00100010_00100010_00100010_00100010_00100010_00011100_00000000;  // O
			7: glyph = 64'b00011110_00100010_00100010_00011110_00100010_00100010_00011110_00000000;  // B
			8: glyph = 64'b00011100_00100010_00100010_00100010_00100010_00100010_00100010_00000000;  // U
			9: glyph = 64'b00111110_00001000_00001000_00001000_00001000_00001000_00111110_00000000;  // I
			10:glyph = 64'b00011100_00100010_00000010_00000010_00000010_00100010_00011100_00000000;  // C
			12:glyph = 64'b00000000_00011000_00011000_00000000_00000000_00011000_00011000_00000000;  // Colon
			
			// Number Glyphs
			13:glyph = 64'b00011100_00100010_00100010_00101010_00100010_00100010_00011100_00000000;  // 0 
			14:glyph = 64'b01111100_00010000_00010000_00010000_00010100_00011000_00010000_00000000;  // 1
			15:glyph = 64'b00111110_00000100_00001000_00010000_00100010_00100010_00011100_00000000;  // 2 
			16:glyph = 64'b00011100_00100010_00100000_00011100_00100000_00100010_00011100_00000000;  // 3
			17:glyph = 64'b00100000_00100000_00100000_00111100_00100100_00100100_00100100_00000000;  // 4 
			18:glyph = 64'b00011110_00100000_00100000_00011110_00000010_00000010_00111110_00000000;  // 5 
			19:glyph = 64'b00011100_00100010_00100010_00011110_00000010_00000100_00111000_00000000;  // 6 
			20:glyph = 64'b00001000_00001000_00001000_00010000_00010000_00100000_00111110_00000000;  // 7
			21:glyph = 64'b00011100_00100010_00100010_00011100_00100010_00100010_00011100_00000000;  // 8 
			22:glyph = 64'b00011100_00100010_00100000_00111100_00100010_00100010_00011100_00000000;  // 9 
			
			// Color Glyphs
			30:glyph = 64'b11111111_11111111_11111111_11111111_11111111_11111111_11111111_11111111;  // White
			31: glyph = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; //Black
			default: glyph = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000; //Black (Should never happen)
		endcase
	
	// Compute the pixel value based on the glyph, row, and column
   // If char_index < 31, extract the bit at the corresponding row and column from the glyph
   // If char_index is 10 (special case), always output 1 (e.g., for a placeholder)
	assign pixel = (char_index < 31) ? glyph[(glyph_row * 8) + glyph_column] : 
	(char_index == 10) ? 1'b1 : 
	1'b0; // Default to 0 for other cases

endmodule